package voq_pkg;

    parameter int VOQ_DEPTH = 8;

endpackage
