`timescale 1ns/1ps

package switch_pkg;

    parameter int NUM_PORTS = 4;

endpackage
