module tx_mac_control #(
    parameter ADDR_W = 6,
    parameter BLOCK_BYTES = 64
)(
    // GMII interface
    output logic gmii_tx_clk_o,
    output logic [DATA_WIDTH-1:0] gmii_tx_data_o,
    output logic gmii_tx_en_o,
    output logic gmii_tx_er_o,
    
    // switch's clk domain
    input logic switch_clk, switch_rst_n,
    
    // mem read ctrl interface
    output logic mem_re_o, mem_start_o,
    output logic [ADDR_W-1:0] mem_start_addr_o,
    input logic [BLOCK_BYTES-1:0][DATA_WIDTH-1:0] frame_data_i, // input data one block at a time
    input logic frame_valid_i, // high for every cycle data is valid
    input logic frame_end_i, // high on last block of frame

    // VOQ signals
    input logic voq_valid_i, // indicates VOQ has valid start ptr
    input logic [ADDR_W-1:0] voq_ptr_i, // starting mem ptr for frame
    output logic voq_ready_o // always high when ready to start frame
);

import rx_tx_pkg::*;
import voq_pkg::*;

// status and debug signals (simulation only)
logic [31:0] tx_frame_count; // # of frames transmitted
logic [31:0] mem_stall_count; // # of times mem read ctrl stalled
logic [31:0] fifo_overflow_count; // # of times FIFO full - switch clk domain
logic [31:0] fifo_underflow_count; // # of times FIFO empty - gmii clk domain

// generate gmii clk
clk_div #(
    .DIVIDE(3) // 3 + 1 = 4, 125MHz from 500MHz switch clk
) gmii_clk_gen (
    .clk_in(switch_clk),
    .rst_n(switch_rst_n),
    .clk_out(gmii_tx_clk_o)
);

// FIFO signals for CDC (switch clk -> GMII)
logic [DATA_WIDTH-1:0] fifo_din; // continous only 
logic fifo_wr_en;
logic fifo_full; logic fifo_empty;
logic fifo_rd_en;

// sync switch clk reset to gmii/PHY clk
logic sync_switch_rst_n;
synchronizer sync_rst(gmii_tx_clk_o, switch_rst_n, sync_switch_rst_n);

// CDC FIFO instance (async FIFO)
async_fifo cdc_fifo (
    .wclk(switch_clk),
    .wrst_n(switch_rst_n),
    .w_en(fifo_wr_en),
    .w_data(fifo_din),
    .w_full(fifo_full),
    
    .rclk(gmii_tx_clk_o),
    .rrst_n(sync_switch_rst_n),
    .r_en(fifo_rd_en),
    .r_data(gmii_tx_data_o),
    .r_empty(fifo_empty)
);

// state machine (switch clk domain) - handles all frame processing
typedef enum logic [1:0] {IDLE, PREAMBLE, DATA, IFG} state_t;

state_t current_state, next_state;

logic [2:0] preamble_ctr, next_preamble_ctr; // 8 bytes
logic [3:0] IFG_ctr, next_IFG_ctr; // 12 bytes
logic [5:0] block_ctr, next_block_ctr; // 64 bytes

// logic should be combinational to avoid cycle delay
// logic next_mem_re_o, next_mem_start_o; 
// logic [ADDR_W-1:0] next_mem_start_addr_o;
// logic next_voq_ready_o;

logic mem_req_flag, next_mem_req_flag; // flag for one cycle mem_re_o
logic prev_mem_re_o; // previous cycle request
logic saved_frame_end_i, next_saved_frame_end_i; // latch frame_end_i when requesting next block
logic mem_stalled; assign mem_stalled = prev_mem_re_o && !frame_valid_i; // mem read requested but no valid data
logic [ADDR_W-1:0] saved_mem_start_addr_o, next_saved_mem_start_addr_o;

// block buffer
logic [BLOCK_BYTES-1:0][DATA_WIDTH-1:0] block_buffer, next_block_buffer;

// status and debug signals
logic [31:0] next_tx_frame_count, next_mem_stall_count;

// // error can be generated by mem stalling during frame transmission or if FIFO underflows during transmission
// logic frame_tx_error, next_frame_tx_error;
// logic [1:0] gmii_tx_error_ff; // sync error to gmii clk domain

always_comb begin
    // default values
    next_state = current_state;
    next_preamble_ctr = preamble_ctr;
    next_IFG_ctr = IFG_ctr;
    next_block_ctr = block_ctr;
    fifo_wr_en = 1'b0;
    mem_re_o = 1'b0;
    mem_start_o = 1'b0;
    mem_start_addr_o = 0;
    voq_ready_o = 1'b0;
    next_saved_mem_start_addr_o = saved_mem_start_addr_o;
    next_block_buffer = block_buffer;
    next_mem_req_flag = mem_req_flag;
    // next_frame_tx_error = 1'b0;
    next_saved_frame_end_i = saved_frame_end_i;
    next_tx_frame_count = tx_frame_count;
    next_mem_stall_count = mem_stall_count;
    fifo_din = 0; // default data

    case (current_state)
        IDLE: begin
            if (!voq_valid_i && (block_ctr == 1)) voq_ready_o = 1'b1; // tell voq ready for next frame
            else begin
                if (block_ctr == 1) begin // use block_ctr == 1 as flag that req has not been sent yet
                    $display("TX MAC CTRL: Starting frame transmission from VOQ ptr 0x%0h", voq_ptr_i);
                    mem_start_addr_o = voq_ptr_i; // feed voq starting addr to mem read ctrl
                    next_saved_mem_start_addr_o = voq_ptr_i; // save starting addr
                    mem_start_o = 1'b1; // start signal
                    mem_re_o = 1'b1; 
                    next_block_ctr = 0; // indicate req has been sent
                end else begin
                    if (mem_stalled) begin // mem is stalled, wait in IDLE instead of jumping to preamble early
                        $display("TX MAC CTRL: Memory read stalled while starting frame transmission, mem_stalled = pre_mem_re_o = %b && !frame_valid_i = %b", prev_mem_re_o, !frame_valid_i);
                        mem_start_addr_o = saved_mem_start_addr_o;
                        mem_start_o = 1'b1; // keep start high too
                        mem_re_o = 1'b1; 
                        next_mem_stall_count = mem_stall_count + 1;
                    end else begin // mem ready, jump to preamble
                        $display("TX MAC CTRL: Memory read ready, beginning frame transmission");
                        next_block_buffer = frame_data_i;
                        next_saved_frame_end_i = frame_end_i; // set frame_end_i for first cycle

                        fifo_din = PREAMBLE_BYTE; // immediately begin sending preamble
                        fifo_wr_en = 1'b1;
                        next_preamble_ctr = 1; // reset ctr

                        next_state = PREAMBLE;
                    end
                end
            end
        end
        PREAMBLE: begin // write 7 preamble bytes + 1 SFD byte
            // latch entire block on first cycle

            if (!fifo_full) begin
                if (preamble_ctr < 7) begin 
                    fifo_din = PREAMBLE_BYTE;
                    $display("TX MAC CTRL: Sending preamble byte at preamble_ctr %0d", preamble_ctr);
                end else begin
                    fifo_din = SFD_BYTE;
                    next_state = DATA;
                    $display("TX MAC CTRL: Sending SFD byte at preamble_ctr %0d", preamble_ctr);
                end
                fifo_wr_en = 1'b1;
                next_preamble_ctr = preamble_ctr + 1;
            end
        end
        DATA: begin // frame_data_i[63] is the footer byte, ignore
            if ((block_ctr == 61) && !saved_frame_end_i) begin // request next block if not last block
                if (!mem_req_flag) begin 
                    mem_re_o = 1'b1; // only assert mem_re_o for one cycle
                    next_saved_frame_end_i = frame_end_i; // latch current frame_end_i before it's updated
                    next_mem_req_flag = 1'b1;
                end else if (mem_stalled) begin 
                    mem_re_o = 1'b1; // stuck here for multiple cycles, so only keep asserting mem_re_o if stalled
                    next_saved_frame_end_i = frame_end_i; // latch current frame_end_i before it's updated
                end
            end else if (block_ctr == 62) begin
                next_mem_req_flag = 1'b0; // reset mem req flag
                if (saved_frame_end_i && !fifo_full) begin // finish writing last byte, then move to IFG
                    next_tx_frame_count = tx_frame_count + 1;
                    next_state = IFG;
                end else if (mem_stalled) begin // mem stalled, stay and don't reset block_ctr 
                    mem_re_o = 1'b1; 
                    next_mem_stall_count = mem_stall_count + 1;
                end else if (!fifo_full) begin // only latch next block if not last block + mem not stalled + last data has gone out
                    next_block_buffer = frame_data_i; // latch next block
                end
            end 

            if (!fifo_full) begin // only write with new data available + fifo not full, also don't update block ctr unless data written
                fifo_din = block_buffer[block_ctr];
                fifo_wr_en = 1'b1;
                next_block_ctr = block_ctr + 1;
            end
        end
        IFG: begin // maintain 12-byte IFG
            next_IFG_ctr = IFG_ctr + 1;
            if (IFG_ctr == 11) begin // wait 11 times then go to IDLE (total 12 bytes)
                voq_ready_o = 1'b1;
                next_IFG_ctr = 0;
                next_block_ctr = 1; // use 1 as a flag
                next_state = IDLE;
            end
        end
        default: next_state = IDLE;
    endcase
end

// state machine (switch clk domain) - seq logic
always_ff @(posedge switch_clk or negedge switch_rst_n) begin
    if (!switch_rst_n) begin
        current_state <= IDLE;
        // mem_re_o <= 0;
        // mem_start_o <= 0;
        // mem_start_addr_o <= 0;
        // voq_ready_o <= 0;
        preamble_ctr <= 0;
        IFG_ctr <= 0;
        block_ctr <= 1;
        block_buffer <= 0;
        saved_mem_start_addr_o <= 0;
        tx_frame_count <= 0;
        mem_stall_count <= 0;
        mem_req_flag <= 0;
        // frame_tx_error <= 0;

        prev_mem_re_o <= 0;
        saved_frame_end_i <= 0;

        fifo_overflow_count <= 0;
    end else begin
        current_state <= next_state;
        // mem_re_o <= next_mem_re_o;
        // mem_start_o <= next_mem_start_o;
        // mem_start_addr_o <= next_mem_start_addr_o;
        // voq_ready_o <= next_voq_ready_o;
        preamble_ctr <= next_preamble_ctr;
        IFG_ctr <= next_IFG_ctr;
        block_ctr <= next_block_ctr;
        block_buffer <= next_block_buffer;
        saved_mem_start_addr_o <= next_saved_mem_start_addr_o;
        tx_frame_count <= next_tx_frame_count;
        mem_stall_count <= next_mem_stall_count;
        mem_req_flag <= next_mem_req_flag;
        // frame_tx_error <= next_frame_tx_error;

        prev_mem_re_o <= mem_re_o;
        saved_frame_end_i <= next_saved_frame_end_i;
        
        // debug counter
        if (fifo_full) fifo_overflow_count <= fifo_overflow_count + 1;
    end
end

// simple output logic (gmii clk domain) - just read from FIFO and output
logic prev_fifo_rd_en;
assign fifo_rd_en = !fifo_empty; // continuous read when data available
assign gmii_tx_en_o = prev_fifo_rd_en; // tx_en follows
assign gmii_tx_er_o = fifo_empty && !frame_end_i; // error if fifo underflow, could be from mem stalling during frame transmission, assume empty on frame end is ok, if not, rx will catch it with crc error 

// simple gmii
always_ff @(posedge gmii_tx_clk_o or negedge sync_switch_rst_n) begin
    if (!sync_switch_rst_n) begin
        fifo_underflow_count <= 0;
        prev_fifo_rd_en <= 0;
    end else begin
        prev_fifo_rd_en <= fifo_rd_en;

        // gmii_tx_error_ff <= {gmii_tx_error_ff[0], frame_tx_error};

        // debug
        if (fifo_empty) fifo_underflow_count <= fifo_underflow_count + 1;
    end
end

endmodule
